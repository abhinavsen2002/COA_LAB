`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:52:44 10/26/2022 
// Design Name: 
// Module Name:    diff 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module diff(
	input [31:0] a,
	input [31:0] b,
	output reg [31:0] i
    );

	reg [31:0] x;
	always@(*) begin
		x = a ^ b;
		i[0] <= x[0];
		// The mountain below is obviously written via python
		i[1] <= ~x[0] & x[1];
		i[2] <= ~x[0] & ~x[1] & x[2];
		i[3] <= ~x[0] & ~x[1] & ~x[2] & x[3];
		i[4] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & x[4];
		i[5] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & x[5];
		i[6] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & x[6];
		i[7] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & x[7];
		i[8] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & x[8];
		i[9] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & x[9];
		i[10] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & x[10];
		i[11] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & x[11];
		i[12] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & x[12];
		i[13] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & x[13];
		i[14] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & x[14];
		i[15] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & x[15];
		i[16] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & x[16];
		i[17] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & x[17];
		i[18] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & x[18];
		i[19] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & x[19];
		i[20] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & x[20];
		i[21] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & x[21];
		i[22] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & x[22];
		i[23] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & x[23];
		i[24] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & x[24];
		i[25] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & x[25];
		i[26] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & x[26];
		i[27] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & x[27];
		i[28] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & x[28];
		i[29] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & x[29];
		i[30] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & x[30];
		i[31] <= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & x[31];
		
	end
	
endmodule
